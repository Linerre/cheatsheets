`timescale 1ns / 1ps
  module (
     input wire        clk,
     input wire        reset,
     input wire        btn_e,
     input wire        btn_w,
     input wire        btn_s,
     input wire        btn_n,
     output reg [15:0] LED,
     output wire [3:0] ANODE,
     output wire [6:0] CATHODE
  );

     // debounce btn

     // spot btn

     // fsm

     // output
  endmodule
